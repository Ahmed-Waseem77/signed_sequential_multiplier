

`resetall
`timescale 1ns/10ps


module signed_sequential_multiplier_tb;



endmodule