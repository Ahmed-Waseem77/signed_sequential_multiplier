//
// Verilog Module signed_sequential_multiplier_lib.prev_mulr_reg
//
// Created:
//          by - ahmed.UNKNOWN (WES-HPOMEN)
//          at - 18:11:10 04/30/2023
//
// using Mentor Graphics HDL Designer(TM) 2023.1 Built on 19 Jan 2023 at 15:19:29
//

`resetall
`timescale 1ns/10ps
module prev_mulr_reg( 
   // Port Declarations
   input   wire    [7:0]   multiplicand, 
   output  wire    [15:0]  previous_mulr
);


// Internal Declarations




// ### Please start your Verilog code here ### 

endmodule
